##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Sun Apr 18 01:54:53 2021
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO aesbuffer
  CLASS BLOCK ;
  SIZE 168.150000 BY 167.720000 ;
  FOREIGN aesbuffer 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.880000 167.650000 52.950000 167.720000 ;
    END
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.930000 167.650000 52.000000 167.720000 ;
    END
  END resetn
  PIN addr_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 83.280000 167.650000 83.350000 167.720000 ;
    END
  END addr_in[31]
  PIN addr_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.330000 167.650000 82.400000 167.720000 ;
    END
  END addr_in[30]
  PIN addr_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.380000 167.650000 81.450000 167.720000 ;
    END
  END addr_in[29]
  PIN addr_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.430000 167.650000 80.500000 167.720000 ;
    END
  END addr_in[28]
  PIN addr_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.480000 167.650000 79.550000 167.720000 ;
    END
  END addr_in[27]
  PIN addr_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.530000 167.650000 78.600000 167.720000 ;
    END
  END addr_in[26]
  PIN addr_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.580000 167.650000 77.650000 167.720000 ;
    END
  END addr_in[25]
  PIN addr_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.630000 167.650000 76.700000 167.720000 ;
    END
  END addr_in[24]
  PIN addr_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.680000 167.650000 75.750000 167.720000 ;
    END
  END addr_in[23]
  PIN addr_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.730000 167.650000 74.800000 167.720000 ;
    END
  END addr_in[22]
  PIN addr_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.780000 167.650000 73.850000 167.720000 ;
    END
  END addr_in[21]
  PIN addr_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.830000 167.650000 72.900000 167.720000 ;
    END
  END addr_in[20]
  PIN addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 71.880000 167.650000 71.950000 167.720000 ;
    END
  END addr_in[19]
  PIN addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.930000 167.650000 71.000000 167.720000 ;
    END
  END addr_in[18]
  PIN addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.980000 167.650000 70.050000 167.720000 ;
    END
  END addr_in[17]
  PIN addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.030000 167.650000 69.100000 167.720000 ;
    END
  END addr_in[16]
  PIN addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.080000 167.650000 68.150000 167.720000 ;
    END
  END addr_in[15]
  PIN addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.130000 167.650000 67.200000 167.720000 ;
    END
  END addr_in[14]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.180000 167.650000 66.250000 167.720000 ;
    END
  END addr_in[13]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.230000 167.650000 65.300000 167.720000 ;
    END
  END addr_in[12]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.280000 167.650000 64.350000 167.720000 ;
    END
  END addr_in[11]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.330000 167.650000 63.400000 167.720000 ;
    END
  END addr_in[10]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.380000 167.650000 62.450000 167.720000 ;
    END
  END addr_in[9]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.430000 167.650000 61.500000 167.720000 ;
    END
  END addr_in[8]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.480000 167.650000 60.550000 167.720000 ;
    END
  END addr_in[7]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.530000 167.650000 59.600000 167.720000 ;
    END
  END addr_in[6]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.580000 167.650000 58.650000 167.720000 ;
    END
  END addr_in[5]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.630000 167.650000 57.700000 167.720000 ;
    END
  END addr_in[4]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.680000 167.650000 56.750000 167.720000 ;
    END
  END addr_in[3]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.730000 167.650000 55.800000 167.720000 ;
    END
  END addr_in[2]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.780000 167.650000 54.850000 167.720000 ;
    END
  END addr_in[1]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.830000 167.650000 53.900000 167.720000 ;
    END
  END addr_in[0]
  PIN mr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.230000 167.650000 84.300000 167.720000 ;
    END
  END mr
  PIN mw
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.180000 167.650000 85.250000 167.720000 ;
    END
  END mw
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.580000 167.650000 115.650000 167.720000 ;
    END
  END data_in[31]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 114.630000 167.650000 114.700000 167.720000 ;
    END
  END data_in[30]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.680000 167.650000 113.750000 167.720000 ;
    END
  END data_in[29]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 112.730000 167.650000 112.800000 167.720000 ;
    END
  END data_in[28]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.780000 167.650000 111.850000 167.720000 ;
    END
  END data_in[27]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.830000 167.650000 110.900000 167.720000 ;
    END
  END data_in[26]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.880000 167.650000 109.950000 167.720000 ;
    END
  END data_in[25]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.930000 167.650000 109.000000 167.720000 ;
    END
  END data_in[24]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.980000 167.650000 108.050000 167.720000 ;
    END
  END data_in[23]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.030000 167.650000 107.100000 167.720000 ;
    END
  END data_in[22]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.080000 167.650000 106.150000 167.720000 ;
    END
  END data_in[21]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.130000 167.650000 105.200000 167.720000 ;
    END
  END data_in[20]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.180000 167.650000 104.250000 167.720000 ;
    END
  END data_in[19]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.230000 167.650000 103.300000 167.720000 ;
    END
  END data_in[18]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.280000 167.650000 102.350000 167.720000 ;
    END
  END data_in[17]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.330000 167.650000 101.400000 167.720000 ;
    END
  END data_in[16]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.380000 167.650000 100.450000 167.720000 ;
    END
  END data_in[15]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.430000 167.650000 99.500000 167.720000 ;
    END
  END data_in[14]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.480000 167.650000 98.550000 167.720000 ;
    END
  END data_in[13]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.530000 167.650000 97.600000 167.720000 ;
    END
  END data_in[12]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.580000 167.650000 96.650000 167.720000 ;
    END
  END data_in[11]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.630000 167.650000 95.700000 167.720000 ;
    END
  END data_in[10]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.680000 167.650000 94.750000 167.720000 ;
    END
  END data_in[9]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.730000 167.650000 93.800000 167.720000 ;
    END
  END data_in[8]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.780000 167.650000 92.850000 167.720000 ;
    END
  END data_in[7]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.830000 167.650000 91.900000 167.720000 ;
    END
  END data_in[6]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.880000 167.650000 90.950000 167.720000 ;
    END
  END data_in[5]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.930000 167.650000 90.000000 167.720000 ;
    END
  END data_in[4]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.980000 167.650000 89.050000 167.720000 ;
    END
  END data_in[3]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.030000 167.650000 88.100000 167.720000 ;
    END
  END data_in[2]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.080000 167.650000 87.150000 167.720000 ;
    END
  END data_in[1]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.130000 167.650000 86.200000 167.720000 ;
    END
  END data_in[0]
  PIN data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 62.195000 168.150000 62.265000 ;
    END
  END data_out[31]
  PIN data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 63.595000 168.150000 63.665000 ;
    END
  END data_out[30]
  PIN data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 64.995000 168.150000 65.065000 ;
    END
  END data_out[29]
  PIN data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 66.395000 168.150000 66.465000 ;
    END
  END data_out[28]
  PIN data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 67.795000 168.150000 67.865000 ;
    END
  END data_out[27]
  PIN data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 69.195000 168.150000 69.265000 ;
    END
  END data_out[26]
  PIN data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 70.595000 168.150000 70.665000 ;
    END
  END data_out[25]
  PIN data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 71.995000 168.150000 72.065000 ;
    END
  END data_out[24]
  PIN data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 73.395000 168.150000 73.465000 ;
    END
  END data_out[23]
  PIN data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 74.795000 168.150000 74.865000 ;
    END
  END data_out[22]
  PIN data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 76.195000 168.150000 76.265000 ;
    END
  END data_out[21]
  PIN data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 77.595000 168.150000 77.665000 ;
    END
  END data_out[20]
  PIN data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 78.995000 168.150000 79.065000 ;
    END
  END data_out[19]
  PIN data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 80.395000 168.150000 80.465000 ;
    END
  END data_out[18]
  PIN data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 81.795000 168.150000 81.865000 ;
    END
  END data_out[17]
  PIN data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 83.195000 168.150000 83.265000 ;
    END
  END data_out[16]
  PIN data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 84.595000 168.150000 84.665000 ;
    END
  END data_out[15]
  PIN data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 85.995000 168.150000 86.065000 ;
    END
  END data_out[14]
  PIN data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 87.395000 168.150000 87.465000 ;
    END
  END data_out[13]
  PIN data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 88.795000 168.150000 88.865000 ;
    END
  END data_out[12]
  PIN data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 90.195000 168.150000 90.265000 ;
    END
  END data_out[11]
  PIN data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 91.595000 168.150000 91.665000 ;
    END
  END data_out[10]
  PIN data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 92.995000 168.150000 93.065000 ;
    END
  END data_out[9]
  PIN data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 94.395000 168.150000 94.465000 ;
    END
  END data_out[8]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 95.795000 168.150000 95.865000 ;
    END
  END data_out[7]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 97.195000 168.150000 97.265000 ;
    END
  END data_out[6]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 98.595000 168.150000 98.665000 ;
    END
  END data_out[5]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 99.995000 168.150000 100.065000 ;
    END
  END data_out[4]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 101.395000 168.150000 101.465000 ;
    END
  END data_out[3]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 102.795000 168.150000 102.865000 ;
    END
  END data_out[2]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 104.195000 168.150000 104.265000 ;
    END
  END data_out[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.080000 105.595000 168.150000 105.665000 ;
    END
  END data_out[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal2 ;
      RECT 115.720000 167.580000 168.150000 167.720000 ;
      RECT 114.770000 167.580000 115.510000 167.720000 ;
      RECT 113.820000 167.580000 114.560000 167.720000 ;
      RECT 112.870000 167.580000 113.610000 167.720000 ;
      RECT 111.920000 167.580000 112.660000 167.720000 ;
      RECT 110.970000 167.580000 111.710000 167.720000 ;
      RECT 110.020000 167.580000 110.760000 167.720000 ;
      RECT 109.070000 167.580000 109.810000 167.720000 ;
      RECT 108.120000 167.580000 108.860000 167.720000 ;
      RECT 107.170000 167.580000 107.910000 167.720000 ;
      RECT 106.220000 167.580000 106.960000 167.720000 ;
      RECT 105.270000 167.580000 106.010000 167.720000 ;
      RECT 104.320000 167.580000 105.060000 167.720000 ;
      RECT 103.370000 167.580000 104.110000 167.720000 ;
      RECT 102.420000 167.580000 103.160000 167.720000 ;
      RECT 101.470000 167.580000 102.210000 167.720000 ;
      RECT 100.520000 167.580000 101.260000 167.720000 ;
      RECT 99.570000 167.580000 100.310000 167.720000 ;
      RECT 98.620000 167.580000 99.360000 167.720000 ;
      RECT 97.670000 167.580000 98.410000 167.720000 ;
      RECT 96.720000 167.580000 97.460000 167.720000 ;
      RECT 95.770000 167.580000 96.510000 167.720000 ;
      RECT 94.820000 167.580000 95.560000 167.720000 ;
      RECT 93.870000 167.580000 94.610000 167.720000 ;
      RECT 92.920000 167.580000 93.660000 167.720000 ;
      RECT 91.970000 167.580000 92.710000 167.720000 ;
      RECT 91.020000 167.580000 91.760000 167.720000 ;
      RECT 90.070000 167.580000 90.810000 167.720000 ;
      RECT 89.120000 167.580000 89.860000 167.720000 ;
      RECT 88.170000 167.580000 88.910000 167.720000 ;
      RECT 87.220000 167.580000 87.960000 167.720000 ;
      RECT 86.270000 167.580000 87.010000 167.720000 ;
      RECT 85.320000 167.580000 86.060000 167.720000 ;
      RECT 84.370000 167.580000 85.110000 167.720000 ;
      RECT 83.420000 167.580000 84.160000 167.720000 ;
      RECT 82.470000 167.580000 83.210000 167.720000 ;
      RECT 81.520000 167.580000 82.260000 167.720000 ;
      RECT 80.570000 167.580000 81.310000 167.720000 ;
      RECT 79.620000 167.580000 80.360000 167.720000 ;
      RECT 78.670000 167.580000 79.410000 167.720000 ;
      RECT 77.720000 167.580000 78.460000 167.720000 ;
      RECT 76.770000 167.580000 77.510000 167.720000 ;
      RECT 75.820000 167.580000 76.560000 167.720000 ;
      RECT 74.870000 167.580000 75.610000 167.720000 ;
      RECT 73.920000 167.580000 74.660000 167.720000 ;
      RECT 72.970000 167.580000 73.710000 167.720000 ;
      RECT 72.020000 167.580000 72.760000 167.720000 ;
      RECT 71.070000 167.580000 71.810000 167.720000 ;
      RECT 70.120000 167.580000 70.860000 167.720000 ;
      RECT 69.170000 167.580000 69.910000 167.720000 ;
      RECT 68.220000 167.580000 68.960000 167.720000 ;
      RECT 67.270000 167.580000 68.010000 167.720000 ;
      RECT 66.320000 167.580000 67.060000 167.720000 ;
      RECT 65.370000 167.580000 66.110000 167.720000 ;
      RECT 64.420000 167.580000 65.160000 167.720000 ;
      RECT 63.470000 167.580000 64.210000 167.720000 ;
      RECT 62.520000 167.580000 63.260000 167.720000 ;
      RECT 61.570000 167.580000 62.310000 167.720000 ;
      RECT 60.620000 167.580000 61.360000 167.720000 ;
      RECT 59.670000 167.580000 60.410000 167.720000 ;
      RECT 58.720000 167.580000 59.460000 167.720000 ;
      RECT 57.770000 167.580000 58.510000 167.720000 ;
      RECT 56.820000 167.580000 57.560000 167.720000 ;
      RECT 55.870000 167.580000 56.610000 167.720000 ;
      RECT 54.920000 167.580000 55.660000 167.720000 ;
      RECT 53.970000 167.580000 54.710000 167.720000 ;
      RECT 53.020000 167.580000 53.760000 167.720000 ;
      RECT 52.070000 167.580000 52.810000 167.720000 ;
      RECT 0.000000 167.580000 51.860000 167.720000 ;
      RECT 0.000000 105.735000 168.150000 167.580000 ;
      RECT 0.000000 105.525000 168.010000 105.735000 ;
      RECT 0.000000 104.335000 168.150000 105.525000 ;
      RECT 0.000000 104.125000 168.010000 104.335000 ;
      RECT 0.000000 102.935000 168.150000 104.125000 ;
      RECT 0.000000 102.725000 168.010000 102.935000 ;
      RECT 0.000000 101.535000 168.150000 102.725000 ;
      RECT 0.000000 101.325000 168.010000 101.535000 ;
      RECT 0.000000 100.135000 168.150000 101.325000 ;
      RECT 0.000000 99.925000 168.010000 100.135000 ;
      RECT 0.000000 98.735000 168.150000 99.925000 ;
      RECT 0.000000 98.525000 168.010000 98.735000 ;
      RECT 0.000000 97.335000 168.150000 98.525000 ;
      RECT 0.000000 97.125000 168.010000 97.335000 ;
      RECT 0.000000 95.935000 168.150000 97.125000 ;
      RECT 0.000000 95.725000 168.010000 95.935000 ;
      RECT 0.000000 94.535000 168.150000 95.725000 ;
      RECT 0.000000 94.325000 168.010000 94.535000 ;
      RECT 0.000000 93.135000 168.150000 94.325000 ;
      RECT 0.000000 92.925000 168.010000 93.135000 ;
      RECT 0.000000 91.735000 168.150000 92.925000 ;
      RECT 0.000000 91.525000 168.010000 91.735000 ;
      RECT 0.000000 90.335000 168.150000 91.525000 ;
      RECT 0.000000 90.125000 168.010000 90.335000 ;
      RECT 0.000000 88.935000 168.150000 90.125000 ;
      RECT 0.000000 88.725000 168.010000 88.935000 ;
      RECT 0.000000 87.535000 168.150000 88.725000 ;
      RECT 0.000000 87.325000 168.010000 87.535000 ;
      RECT 0.000000 86.135000 168.150000 87.325000 ;
      RECT 0.000000 85.925000 168.010000 86.135000 ;
      RECT 0.000000 84.735000 168.150000 85.925000 ;
      RECT 0.000000 84.525000 168.010000 84.735000 ;
      RECT 0.000000 83.335000 168.150000 84.525000 ;
      RECT 0.000000 83.125000 168.010000 83.335000 ;
      RECT 0.000000 81.935000 168.150000 83.125000 ;
      RECT 0.000000 81.725000 168.010000 81.935000 ;
      RECT 0.000000 80.535000 168.150000 81.725000 ;
      RECT 0.000000 80.325000 168.010000 80.535000 ;
      RECT 0.000000 79.135000 168.150000 80.325000 ;
      RECT 0.000000 78.925000 168.010000 79.135000 ;
      RECT 0.000000 77.735000 168.150000 78.925000 ;
      RECT 0.000000 77.525000 168.010000 77.735000 ;
      RECT 0.000000 76.335000 168.150000 77.525000 ;
      RECT 0.000000 76.125000 168.010000 76.335000 ;
      RECT 0.000000 74.935000 168.150000 76.125000 ;
      RECT 0.000000 74.725000 168.010000 74.935000 ;
      RECT 0.000000 73.535000 168.150000 74.725000 ;
      RECT 0.000000 73.325000 168.010000 73.535000 ;
      RECT 0.000000 72.135000 168.150000 73.325000 ;
      RECT 0.000000 71.925000 168.010000 72.135000 ;
      RECT 0.000000 70.735000 168.150000 71.925000 ;
      RECT 0.000000 70.525000 168.010000 70.735000 ;
      RECT 0.000000 69.335000 168.150000 70.525000 ;
      RECT 0.000000 69.125000 168.010000 69.335000 ;
      RECT 0.000000 67.935000 168.150000 69.125000 ;
      RECT 0.000000 67.725000 168.010000 67.935000 ;
      RECT 0.000000 66.535000 168.150000 67.725000 ;
      RECT 0.000000 66.325000 168.010000 66.535000 ;
      RECT 0.000000 65.135000 168.150000 66.325000 ;
      RECT 0.000000 64.925000 168.010000 65.135000 ;
      RECT 0.000000 63.735000 168.150000 64.925000 ;
      RECT 0.000000 63.525000 168.010000 63.735000 ;
      RECT 0.000000 62.335000 168.150000 63.525000 ;
      RECT 0.000000 62.125000 168.010000 62.335000 ;
      RECT 0.000000 0.000000 168.150000 62.125000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 168.150000 167.720000 ;
  END
END aesbuffer

END LIBRARY
